
module	FPGACore
		(
			
		)
	
	always_comb
	begin
	
	end
endmodule 
